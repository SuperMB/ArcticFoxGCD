/*
Copyright (c) 2022, Icii Technologies LLC
All rights reserved.

This source code is licensed under the BSD-style license found in the
LICENSE file in the root directory of this source tree. 
*/

module Registers(      
);





//[CommandReg]
wire [15:0] gcd1;
// [CommandReg]
wire [15:0] gcd2;

//[CommandPulseReg -command StartGCD]
reg startGCD;



                

endmodule
